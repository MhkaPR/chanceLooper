module chanceLooper (
    input clk,
    
);
    
endmodule